`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////


module OR_Gate(a,b,Y);
input wire a,b;
output Y;
assign Y=a|b;
endmodule
