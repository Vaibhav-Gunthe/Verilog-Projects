`timescale 1ns / 1ps


module Mux2x1(
input I0,
input I1,
input Sel,
output Y
    );
    assign Y=Sel ? I0 : I1;
endmodule
