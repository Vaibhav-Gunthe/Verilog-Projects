`timescale 1ns / 1ps

module XOR_Gate(
input a,b,
output wire Y
    );
    assign Y=a^b;
endmodule
